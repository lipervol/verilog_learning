library verilog;
use verilog.vl_types.all;
entity steppluse_vlg_tst is
end steppluse_vlg_tst;
