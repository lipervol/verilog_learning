library verilog;
use verilog.vl_types.all;
entity myname_vlg_tst is
end myname_vlg_tst;
